entity m9_barrel32 is
port (x   : in std_logic_vector(31 downto 0);
      pos : in std_logic_vector( 4 downto 0);
      lnr : in std_logic;
      y   : in end m9_barrel32;
end m9_barrel32;
