type fix824 is array(31 downto 0) of std_logic_vector(31 downto 0);
constant rom_arctan: fix824:= (
  "00000000000000000000000000011111",
  "00000000000000000000000000111111",
  ...
  "00000000000000000000000001111111");
