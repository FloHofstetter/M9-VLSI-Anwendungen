entity m9_artan_rom is
  port (i : in  std_logic_vector(4 downto 0);
        d : out std_logic_vector(31 downto 0));
end m9_artan_rom;
