entity m9_addsub32 is
    port (a, b : in std_logic_vector(31 downto 0);
          ans  : in std_logic;
          y    : in std_logic_vector(31 downto 0));
end m9_barrel;
