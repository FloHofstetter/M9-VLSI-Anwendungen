library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity m9_artan_rom is
  port(i : in  std_logic_vector(4 downto 0);
       d : out std_logic_vector(31 downto 0));
end m9_artan_rom;

architecture Behavioral of m9_artan_rom is
  type fix824 is array(0 to 31) of std_logic_vector(31 downto 0);
  constant rom_arctan: fix824:= (
    x"00_C9_0F_DB",  -- 00 -> 0,785398
    x"00_76_B1_9C",  -- 01 -> 0.463648
    x"00_3E_B6_EC",  -- 02 -> ...
    x"00_1E_D5_BB",  -- 03 -> ...
    x"00_0E_EA_AE",  -- 04 -> ...
    x"00_07_EE_55",  -- 05 -> ...
    x"00_03_EE_EB",  -- 06 -> ...
    x"00_01_FF_FD",  -- 07 -> ...
    x"00_01_00_00",  -- 08 -> ...
    x"00_00_80_00",  -- 09 -> ...
    x"00_00_40_00",  -- 10 -> ...
    x"00_00_20_00",  -- 11 -> ...
    x"00_00_10_00",  -- 12 -> ...
    x"00_00_08_00",  -- 13 -> ...
    x"00_00_04_00",  -- 14 -> ...
    x"00_00_02_00",  -- 15 -> 0.000015
    x"00_00_01_00",  -- 16 -> ...
    x"00_00_00_80",  -- 17 -> ...
    x"00_00_00_40",  -- 18 -> ...
    x"00_00_00_20",  -- 19 -> ...
    x"00_00_00_10",  -- 20 -> ...
    x"00_00_00_08",  -- 21 -> ...
    x"00_00_00_04",  -- 22 -> ...
    x"00_00_00_02",  -- 23 -> ...
    x"00_00_00_01",  -- 24 -> ...
    x"00_00_00_00",  -- 25 -> ...
    x"00_00_00_00",  -- 26 -> ...
    x"00_00_00_00",  -- 27 -> ...
    x"00_00_00_00",  -- 28 -> ...
    x"00_00_00_00",  -- 29 -> ...
    x"00_00_00_00",  -- 30 -> 0.93E-9
    x"00_00_00_00"   -- 31 -> 0.46e-9
  );
begin
  with i select d <=
    rom_arctan(0)  when "00000",  -- 00
    rom_arctan(1)  when "00001",  -- 01
    rom_arctan(2)  when "00010",  -- 02
    rom_arctan(3)  when "00011",  -- 03
    rom_arctan(4)  when "00100",  -- 04
    rom_arctan(5)  when "00101",  -- 05
    rom_arctan(6)  when "00110",  -- 06
    rom_arctan(7)  when "00111",  -- 07
    rom_arctan(8)  when "01000",  -- 08
    rom_arctan(9)  when "01001",  -- 09
    rom_arctan(10) when "01010",  -- 10
    rom_arctan(11) when "01011",  -- 11
    rom_arctan(12) when "01100",  -- 12
    rom_arctan(13) when "01101",  -- 13
    rom_arctan(14) when "01110",  -- 14
    rom_arctan(15) when "01111",  -- 15
    rom_arctan(16) when "10000",  -- 16
    rom_arctan(17) when "10001",  -- 17
    rom_arctan(18) when "10010",  -- 18
    rom_arctan(19) when "10011",  -- 19
    rom_arctan(20) when "10100",  -- 20
    rom_arctan(21) when "10101",  -- 21
    rom_arctan(22) when "10110",  -- 22
    rom_arctan(23) when "10111",  -- 23
    rom_arctan(24) when "11000",  -- 24
    rom_arctan(25) when "11001",  -- 25
    rom_arctan(26) when "11010",  -- 26
    rom_arctan(27) when "11011",  -- 27
    rom_arctan(28) when "11100",  -- 28
    rom_arctan(29) when "11101",  -- 29
    rom_arctan(30) when "11110",  -- 30
    rom_arctan(31) when "11111",  -- 31
  x"00_00_00_00" when others;
end Behavioral;
